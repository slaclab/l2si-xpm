xpm_sim.vhd.axil