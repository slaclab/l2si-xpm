
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;

library surf;
use surf.StdRtlPkg.all;

package FpgaTypePkg is

  constant CPSW_TARBALL_ADDR_C : slv(31 downto 0) := (others=>'0');
  
end FpgaTypePkg;
